module vga(input clk, output hsync, output vsync);
endmodule
